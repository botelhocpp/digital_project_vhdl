LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY sync IS
	PORT(clk: IN STD_LOGIC;
	     a : IN STD_LOGIC;
	     b: OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE rtl OF sync IS
	SIGNAL m: STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";	
	BEGIN
		PROCESS(clk) IS
			BEGIN
				IF RISING_EDGE(clk) THEN
					m <= m(0) & a;
				END IF;
		END PROCESS;
		b <= m(1);
END ARCHITECTURE;

